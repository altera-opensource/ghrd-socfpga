
module altera_ace5lite_cache_coherency_translator #(
	parameter F2H_ADDRESS_WIDTH=40,
	localparam F2H_DATA_WIDTH=256
) (
	input wire axi_clock,
	input wire axi_reset,

	input wire [5-1:0] axi4_fpga2hps_awid,
	input wire [F2H_ADDRESS_WIDTH-1:0] axi4_fpga2hps_awaddr,
	input wire [8-1:0] axi4_fpga2hps_awlen,
	input wire [3-1:0] axi4_fpga2hps_awsize,
	input wire [3-1:0] axi4_fpga2hps_arsize,
	input wire [2-1:0] axi4_fpga2hps_awburst,
	input wire [1-1:0] axi4_fpga2hps_awlock,
	input wire [4-1:0] axi4_fpga2hps_awcache,
	input wire [3-1:0] axi4_fpga2hps_awprot,
	input wire [4-1:0] axi4_fpga2hps_awqos,
	input wire [1-1:0] axi4_fpga2hps_awvalid,
	output wire [1-1:0] axi4_fpga2hps_awready,
	input wire [F2H_DATA_WIDTH-1:0] axi4_fpga2hps_wdata,
	input wire [F2H_DATA_WIDTH/8-1:0] axi4_fpga2hps_wstrb,
	input wire [1-1:0] axi4_fpga2hps_wlast,
	input wire [1-1:0] axi4_fpga2hps_wvalid,
	output wire [1-1:0] axi4_fpga2hps_wready,
	output wire [5-1:0] axi4_fpga2hps_bid,
	output wire [2-1:0] axi4_fpga2hps_bresp,
	output wire [1-1:0] axi4_fpga2hps_bvalid,
	input wire [1-1:0] axi4_fpga2hps_bready,
	input wire [5-1:0] axi4_fpga2hps_arid,
	input wire [F2H_ADDRESS_WIDTH-1:0] axi4_fpga2hps_araddr,
	input wire [8-1:0] axi4_fpga2hps_arlen,
	input wire [2-1:0] axi4_fpga2hps_arburst,
	input wire [1-1:0] axi4_fpga2hps_arlock,
	input wire [4-1:0] axi4_fpga2hps_arcache,
	input wire [3-1:0] axi4_fpga2hps_arprot,
	input wire [4-1:0] axi4_fpga2hps_arqos,
	input wire [1-1:0] axi4_fpga2hps_arvalid,
	output wire [1-1:0] axi4_fpga2hps_arready,
	output wire [5-1:0] axi4_fpga2hps_rid,
	output wire [F2H_DATA_WIDTH-1:0] axi4_fpga2hps_rdata,
	output wire [2-1:0] axi4_fpga2hps_rresp,
	output wire [1-1:0] axi4_fpga2hps_rlast,
	output wire [1-1:0] axi4_fpga2hps_rvalid,
	input wire [1-1:0] axi4_fpga2hps_rready,
	input wire [8-1:0] axi4_fpga2hps_aruser,
	input wire [8-1:0] axi4_fpga2hps_awuser,
	input wire [4-1:0] axi4_fpga2hps_arregion,
	input wire [4-1:0] axi4_fpga2hps_awregion,
	input wire [8-1:0] axi4_fpga2hps_wuser,
	output wire [8-1:0] axi4_fpga2hps_buser,
	output wire [8-1:0] axi4_fpga2hps_ruser,

	output wire [5-1:0] ace5_fpga2hps_awid,
	output wire [F2H_ADDRESS_WIDTH-1:0] ace5_fpga2hps_awaddr,
	output wire [2-1:0] ace5_fpga2hps_awdomain,
	output wire [4-1:0] ace5_fpga2hps_awsnoop,
	output wire [2-1:0] ace5_fpga2hps_awbar,
	output wire [8-1:0] ace5_fpga2hps_awlen,
	output wire [3-1:0] ace5_fpga2hps_awsize,
	output wire [3-1:0] ace5_fpga2hps_arsize,
	output wire [2-1:0] ace5_fpga2hps_awburst,
	output wire [1-1:0] ace5_fpga2hps_awlock,
	output wire [4-1:0] ace5_fpga2hps_awcache,
	output wire [3-1:0] ace5_fpga2hps_awprot,
	output wire [4-1:0] ace5_fpga2hps_awqos,
	output wire [1-1:0] ace5_fpga2hps_awvalid,
	input wire [1-1:0] ace5_fpga2hps_awready,
	output wire [F2H_DATA_WIDTH-1:0] ace5_fpga2hps_wdata,
	output wire [F2H_DATA_WIDTH/8-1:0] ace5_fpga2hps_wstrb,
	output wire [1-1:0] ace5_fpga2hps_wlast,
	output wire [1-1:0] ace5_fpga2hps_wvalid,
	input wire [1-1:0] ace5_fpga2hps_wready,
	output wire [11-1:0] ace5_fpga2hps_awstashnid,
	output wire [1-1:0] ace5_fpga2hps_awstashniden,
	output wire [5-1:0] ace5_fpga2hps_awstashlpid,
	output wire [1-1:0] ace5_fpga2hps_awstashlpiden,
	output wire [6-1:0] ace5_fpga2hps_awatop,
	input wire [5-1:0] ace5_fpga2hps_bid,
	input wire [2-1:0] ace5_fpga2hps_bresp,
	input wire [1-1:0] ace5_fpga2hps_bvalid,
	output wire [1-1:0] ace5_fpga2hps_bready,
	output wire [5-1:0] ace5_fpga2hps_arid,
	output wire [F2H_ADDRESS_WIDTH-1:0] ace5_fpga2hps_araddr,
	output wire [2-1:0] ace5_fpga2hps_ardomain,
	output wire [4-1:0] ace5_fpga2hps_arsnoop,
	output wire [2-1:0] ace5_fpga2hps_arbar,
	output wire [8-1:0] ace5_fpga2hps_arlen,
	output wire [2-1:0] ace5_fpga2hps_arburst,
	output wire [1-1:0] ace5_fpga2hps_arlock,
	output wire [4-1:0] ace5_fpga2hps_arcache,
	output wire [3-1:0] ace5_fpga2hps_arprot,
	output wire [4-1:0] ace5_fpga2hps_arqos,
	output wire [1-1:0] ace5_fpga2hps_arvalid,
	input wire [1-1:0] ace5_fpga2hps_arready,
	input wire [5-1:0] ace5_fpga2hps_rid,
	input wire [F2H_DATA_WIDTH-1:0] ace5_fpga2hps_rdata,
	input wire [2-1:0] ace5_fpga2hps_rresp,
	input wire [1-1:0] ace5_fpga2hps_rlast,
	input wire [1-1:0] ace5_fpga2hps_rvalid,
	output wire [1-1:0] ace5_fpga2hps_rready,
	output wire [8-1:0] ace5_fpga2hps_aruser,
	output wire [8-1:0] ace5_fpga2hps_awuser,
	output wire [4-1:0] ace5_fpga2hps_arregion,
	output wire [4-1:0] ace5_fpga2hps_awregion,
	output wire [8-1:0] ace5_fpga2hps_wuser,
	input wire [8-1:0] ace5_fpga2hps_buser,
	input wire [8-1:0] ace5_fpga2hps_ruser
);

	assign ace5_fpga2hps_awid = axi4_fpga2hps_awid;
	assign ace5_fpga2hps_awaddr = axi4_fpga2hps_awaddr;
	assign ace5_fpga2hps_awdomain = '0;
	assign ace5_fpga2hps_awsnoop = '0;
	assign ace5_fpga2hps_awbar = '0;
	assign ace5_fpga2hps_awlen = axi4_fpga2hps_awlen;
	assign ace5_fpga2hps_awsize = axi4_fpga2hps_awsize;
	assign ace5_fpga2hps_arsize = axi4_fpga2hps_arsize;
	assign ace5_fpga2hps_awburst = axi4_fpga2hps_awburst;
	assign ace5_fpga2hps_awlock = axi4_fpga2hps_awlock;
	assign ace5_fpga2hps_awcache = axi4_fpga2hps_awcache;
	assign ace5_fpga2hps_awprot = axi4_fpga2hps_awprot;
	assign ace5_fpga2hps_awqos = axi4_fpga2hps_awqos;
	assign ace5_fpga2hps_awvalid = axi4_fpga2hps_awvalid;
	assign axi4_fpga2hps_awready = ace5_fpga2hps_awready;
	assign ace5_fpga2hps_wdata = axi4_fpga2hps_wdata;
	assign ace5_fpga2hps_wstrb = axi4_fpga2hps_wstrb;
	assign ace5_fpga2hps_wlast = axi4_fpga2hps_wlast;
	assign ace5_fpga2hps_wvalid = axi4_fpga2hps_wvalid;
	assign axi4_fpga2hps_wready = ace5_fpga2hps_wready;
	assign ace5_fpga2hps_awstashnid = '0;
	assign ace5_fpga2hps_awstashniden = '0;
	assign ace5_fpga2hps_awstashlpid = '0;
	assign ace5_fpga2hps_awstashlpiden = '0;
	assign ace5_fpga2hps_awatop = '0;
	assign axi4_fpga2hps_bid = ace5_fpga2hps_bid;
	assign axi4_fpga2hps_bresp = ace5_fpga2hps_bresp;
	assign axi4_fpga2hps_bvalid = ace5_fpga2hps_bvalid;
	assign ace5_fpga2hps_bready = axi4_fpga2hps_bready;
	assign ace5_fpga2hps_arid = axi4_fpga2hps_arid;
	assign ace5_fpga2hps_araddr = axi4_fpga2hps_araddr;
	assign ace5_fpga2hps_ardomain = '0;
	assign ace5_fpga2hps_arsnoop = '0;
	assign ace5_fpga2hps_arbar = '0;
	assign ace5_fpga2hps_arlen = axi4_fpga2hps_arlen;
	assign ace5_fpga2hps_arburst = axi4_fpga2hps_arburst;
	assign ace5_fpga2hps_arlock = axi4_fpga2hps_arlock;
	assign ace5_fpga2hps_arcache = axi4_fpga2hps_arcache;
	assign ace5_fpga2hps_arprot = axi4_fpga2hps_arprot;
	assign ace5_fpga2hps_arqos = axi4_fpga2hps_arqos;
	assign ace5_fpga2hps_arvalid = axi4_fpga2hps_arvalid;
	assign axi4_fpga2hps_arready = ace5_fpga2hps_arready;
	assign axi4_fpga2hps_rid = ace5_fpga2hps_rid;
	assign axi4_fpga2hps_rdata = ace5_fpga2hps_rdata;
	assign axi4_fpga2hps_rresp = ace5_fpga2hps_rresp;
	assign axi4_fpga2hps_rlast = ace5_fpga2hps_rlast;
	assign axi4_fpga2hps_rvalid = ace5_fpga2hps_rvalid;
	assign ace5_fpga2hps_rready = axi4_fpga2hps_rready;
	assign ace5_fpga2hps_aruser = axi4_fpga2hps_aruser;
	assign ace5_fpga2hps_awuser = axi4_fpga2hps_awuser;
	assign ace5_fpga2hps_arregion = axi4_fpga2hps_arregion;
	assign ace5_fpga2hps_awregion = axi4_fpga2hps_awregion;
	assign ace5_fpga2hps_wuser = axi4_fpga2hps_wuser;
	assign axi4_fpga2hps_buser = ace5_fpga2hps_buser;
	assign axi4_fpga2hps_rdata = ace5_fpga2hps_rdata;
	assign axi4_fpga2hps_ruser = ace5_fpga2hps_ruser;

endmodule;
